interface inf(input bit clk,rst);
  logic wen;
  logic ren;
  logic [3:0] addr;
  logic [7:0] wdata;
  logic [7:0] rdata;
  
  
  
  
endinterface


